`ifndef ENABLE_CONTROLLER_UVC_PKG_SV
`define ENABLE_CONTROLLER_UVC_PKG_SV

package enable_controller_uvc_pkg;


  `include "uvm_macros.svh"
  import uvm_pkg::*;


  `include "enable_controller_uvc_sequence_item.sv"
  `include "enable_controller_uvc_config.sv"
  `include "enable_controller_uvc_sequencer.sv"
  `include "enable_controller_uvc_monitor.sv"
  `include "enable_controller_uvc_driver.sv"
  `include "enable_controller_uvc_agent.sv"



// AGREGAR LIBRERIA
  `include "enable_controller_uvc_sequence_base.sv"

endpackage:enable_controller_uvc_pkg


`endif //ENABLE_CONTROLLER_UVC_PKG_SV